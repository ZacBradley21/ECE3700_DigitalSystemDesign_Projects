`timescale 1ns/1ps
module testbench ();
   
   // DECLARE SIGNALS
   reg clk;     // "reg" type signals are  controlled
   reg signed [7:0] a;  // by the testbench
   reg signed [7:0] b;  // by the testbench

   integer clk_count = 0;   
   
   // INITIAL SIGNAL CONFIGURATION:
   initial begin
      clk = 0;      
      a   = 0;
      b   = 0;
   end

   // GENERATE CLOCK:
   initial forever #10 clk = ~clk;
   
   // CREATE STIMULI:
   always @(posedge clk) begin
      a <= $random();
      b <= $random();
   end

   // WRITE OUTPUT TO CONSOLE:
   integer fid;
   initial fid = $fopen("test_result.txt", "w");
   
   always @(posedge clk) begin
      $write("clk:  %d", clk_count);      
      $write("\ta:  %b", a);
      $write("\tb:  %b", b);
      $write("\n");
      
      $fwrite(fid,"clk:  %d", clk_count);      
      $fwrite(fid,"\ta:  %b", a);
      $fwrite(fid,"\tb:  %b", b);
      $fwrite(fid,"\n");
   end

   // DEFINE WHEN TO TERMINATE SIMULATION:
   always @(posedge clk) begin
      clk_count <= clk_count + 1;
      if (clk_count == 8) begin
	 $fclose(fid);
	 $finish;
      end
   end

   // ADDITIONAL TEST CASES FOR OVERFLOW
   always @(posedge clk) begin
      if (a + b < a || a + b < b) begin
         $display("Overflow occurred on addition: a = %b, a = %d, b = %b, b = %d", a, a, b, b);
      end
      if (b > a) begin
         $display("Overflow occurred on subtraction: a = %b, a = %d, b = %b, b = %d", a, a, b, b);
   end
   end
endmodule // testbench